package shared_pkg;
	  // Correct and error count variables
  integer correct_count=0;
  integer error_count=0;
  logic test_finished;
  parameter FIFO_WIDTH = 16;
parameter FIFO_DEPTH = 8;
endpackage : shared_pkg